
module BoothMultiplier (
    input [31:0] A,
    input [31:0] B,
    output [63:0] F
);

    reg [63:0] product;
    reg [4:0] counter;
    reg [1:0] state;

    // TODO: Implement a 32-bit multiplier using 'Booth's Algorithm'

endmodule
